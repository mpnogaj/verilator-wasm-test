module test();
	logic [7:0] unused_signal;
endmodule